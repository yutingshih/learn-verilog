module Hello;
    initial begin
        $display("Hello world");
        $finish;
    end
endmodule
